`timescale 1ns / 10ps

module tb_booth_multiplier;

  parameter MUL_SIZE = 4;

  reg                          clk;
  reg                          rst_n;
  reg                          start;
  wire                         ready;
  reg                          sign;
  reg signed  [  MUL_SIZE-1:0] a;
  reg signed  [  MUL_SIZE-1:0] b;
  wire signed [2*MUL_SIZE-1:0] y;

  booth_multiplier #(
    .MUL_WIDTH(MUL_SIZE)
  ) mul (
    .clk     (clk),
    .rst_n   (rst_n),
    .start   (start),
    .sign    (sign),
    .data_in1(a),
    .data_in2(b),
    .data_out(y),
    .ready   (ready)
  );

  initial begin
    clk = 1'b0;
    while (1) begin
      clk = ~clk;
      #5;
    end
  end

  initial begin
    start = 'b0;
    rst_n = 'b0;
    #10 rst_n = 'b1;
    #10;

    sign  = 'b0;
    a     = 6;
    b     = 3;
    start = 1'b1;
    #10 start = 1'b0;
    @(posedge ready);
    #10;
    $display("a: %u, b: %u, a*b: %d", $unsigned(a), $unsigned(b), y);
    if (y == ($unsigned(a) * $unsigned(b))) begin
      $display("result successfull");
    end else begin
      $display("wrong result");
    end

    sign  = 'b1;
    a     = -6;
    b     = 3;
    start = 1'b1;
    #10 start = 1'b0;
    @(posedge ready);
    #10;
    $display("a: %d, b: %d, a*b: %d", a, b, y);
    if (y == a * b) begin
      $display("result successfull");
    end else begin
      $display("wrong result");
    end

    sign  = 'b1;
    a     = -6;
    b     = -3;
    start = 1'b1;
    #10 start = 1'b0;
    @(posedge ready);
    #10;
    $display("a: %d, b: %d, a*b: %d", a, b, y);
    if (y == a * b) begin
      $display("result successfull");
    end else begin
      $display("wrong result");
    end

    sign  = 'b1;
    a     = -7;
    b     = -2;
    start = 1'b1;
    #10 start = 1'b0;
    @(posedge ready);
    #10;
    $display("a: %d, b: %d, a*b: %d", a, b, y);
    if (y == a * b) begin
      $display("result successfull");
    end else begin
      $display("wrong result");
    end

    $finish;
  end
endmodule
